`timescale 1ns / 1ps
`default_nettype none

module noDebounce(

    );
endmodule
