
parameter BYTE_SIZE = 8;
parameter ADD = 3'b000;
parameter SLI = 3'b001;
parameter J = 3'b010;
parameter JAL = 3'b011;
parameter LW = 3'b100;
parameter SW = 3'b101;
parameter BEQ = 3'b110;
parameter ADDI = 3'b111;


`define ALU_ADD 3'b000